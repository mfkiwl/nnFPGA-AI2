package mult_core_packege;

    parameter pTYPE_OF_TRANSFORM = "lin"; // other is log


    // mult widths
    parameter ;
    parameter ;
    parameter ;
    parameter ;
    parameter ;

    // adder part 

endpackage