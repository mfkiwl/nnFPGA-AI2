package mult_core_packege;

    // mult widths
    parameter ;
    parameter ;
    parameter ;
    parameter ;
    parameter ;

    // adder part 

endpackage