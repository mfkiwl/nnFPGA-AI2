module mem_model #(
    parameter pIN_DATA_WIDTH = 16 ,
    parameter pMEM_SIZE      = 228
)(
    input                           iclk,
    input [pIN_DATA_WIDTH-1:0]      idata,
    input []
    input []
    input                           ird_en,
    input                           iwr_en,

    output                           odata
);


endmodule