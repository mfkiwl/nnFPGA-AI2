module posit_add_sub #(

)(

);




endmodule 