module top ( 

);

// fsm

// in_mem

// multiply


// out_mem


endmodule 